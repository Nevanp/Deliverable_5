module timing_recovery(
    input clk,
    input signed [17:0] x_in,
    output reg trig
);

endmodule